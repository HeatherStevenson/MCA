BZh91AY&SY�� "߀Ryg���o������`�
�`  h 	LO����A��hh 4 c��4b�` `M0F	��� 0�2h�14�@��`�M4 a��5
?TɓM14�=Bd�h`� ��L�1M00&�#��M @�" 	�14i���O$�$�4b#ڌ
p�(Q�I���KB0L�qa���xrj�,��~�_���}?��>mL���n�x.�?2�m�*-*I5�Z��)&K����.�d������Q�\)��Hܮ04X;��X�3���w�4�3J����d�2�`+**�z���eO��L�f@H$H�$}�[�@ae+t��qd��P��J��hݪ��SJ��tpjrt��-�����v�L��U��o�}�+�.7�E��[�j���6`�bu��bl��=�G~F�ʹq�{	�E%*�O��!�:}��*;:�˭��5�I�ʇ�fc0��fz��H�F����j��_��j�`�Y#bR�Mtj�J�e/|�/ܯ:�j���p��-S��`�jb��I��[�-Km��7>�;N���6�Dnm��x�pHd&o��<O_�yUl��`���]�U'��\� �:_�!�:M�J4(L�-/��,�TU]�hcC#�,��h��J�Q`�	�07�.3 l-��afʻ��K�KL���D��H������|�#���t��v}��-?�M[�Z�m<���36Jk�3����mj�Z��o����u���k&�1t`�����Y�yZlz'�:GoY�c�R�c����bO��2ԅQ��D�.9��w����7�u��H���v�_�q~��Z]�k����uI>v�������oe����ʯ	ɠ��-���j�G�<���me�9f�~�ab�����lE.�l0�ũ�ۧ�����P�����K��/�ߗ���S��k	v2�Tx/�`ʲ�0��0��`,���k�eK���[Z�kz"��g��ZcAn,g{���V�}C�9�}]GQ�b,�s���l2�~[UQN�0d����G?ېô�)��2[�V)-;aQ�Iڍk�R�)�C�;ݔ�G�,�	�����hK�$�g�ه����q���,�Jw1qc'�O�u���wG#��1dr`�'H�z���9��v�8y��V�i�B��1(��[v�,��c�{��+I�U�#�3Fi6���t<�:�`�3���a��'���YIE?YJ�QIqr�xK�ݽS�RIRR/11���;1C��u���P0�9A6��k91GȬI�~q����J,Z3�����yCCMi�J1�/dl߉������B�o���.�������j��kt�߭�w����3��ɹ���_"���>=M�����r�G[��4�=':.���O{{�Ϊ���8�|�G��]�rq9}ʤ�1D~�IP����QH��C�?�x�jf�=�%�f�5�C��d�UI��8T*��K]�1X�W�j�*^���Ʀo;�;�{�k|$���^;�Lo�UU�V���·~"��.-�v't��0ѣ�M$��ٝ�X��ɣS!�������3H׹��>��Qdn�.��Aا����y��le\����t0dm����R�2��}s���t�p��UI:)��JRq��rE8P���