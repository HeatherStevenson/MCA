BZh91AY&SY�T� �_�Py���g߰����P�t%�( ���~����L� �@ `�1 �&	�!��L����&�L�@   �h9�#� �&���0F&D��Ɉh&�i����)�2Ԑ�	V�KD��V�~0lX�_�eB�D�@��5�Y�e/`���F �j�V�L���J�3-y��k�9 ��'-��m� r<Mvԋ%; � �LeΖ.���=�������m=p5�K�!&Gt�91�d	��NԔ��b�Ѕ�;.f�*
0f�&�N�f3,�@E{+&o��-�u�4��� a밌 j�#e�5R�'D6��U6�S]0����F >q(�
9
��$�1B!!�X� ��RG�Z���
!�A��,��9�5(��c���V��I�q�,^YƶӰ�%�ܖ:�3�;�����Sz2v��a�?B��5��V�ȃA�B��L�Q����#򴸄)%i��
f�H�QZJU�J�s���n�Խ��y���
��cС�QXޟ>�����Trb1�p��!n�.���I�HӼM�,� �7�5^)���
�S!A2؎<x��Bz���=��9v��<��s$%�,�Ā���� k� ��;A��ϱ6�2�k��-�\)�ȝ�AC<D0H����(cDj���e��T��Z�%���@@MQhR�p��XӜz�#A��s&s|��s�^Sh{Lɼ��Y!˘�쇼C�һ��� 8$B�x�#�|���,,M*Z4Kڨ2�vC�Tr��O-�r%������-�7���C9��fc:��:F�X��0��YZdNlMr��5:�O��?��`.=�d� ^`�������H�
 �j�`