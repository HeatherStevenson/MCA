BZh91AY&SY�1O� #߀Ryg���o������`�  �    2dшbi���4�&&�h �dɣ��i�0LM4��8ɓF!���`��i�q�&�CL	��14�@j&�j�4hi���M�4 I&�ɐ&��I��m&���<�8b
�(���
%�	&�I8���?7�xt��,~}O�����ߎo����2�4f��ݟ<M�ܴ��eE�I&���/�$�t�B�b�&J)_�S�ڮ�J��H�gm��>W��������|��ܿ����i>��W���glX��K�i�V5����d\����~����l�ދZʳ���{S�|��loº:i�%ZN�e�9��O>;���]Փ��\*��i�dV̸ްa�rߋ=1�N�n
�NǊ�M������OШֲ��1��M�))]\�w�&c$u�m�v�Y��.aW�0���f3	9X��6i'�H�-cZ�*�D��t�VM$��~�[7����?v<��^Ū��#GNn4���k�M/�q�n�������r�S��x���UM�R��UUJ����Yu-=������]+m�3�^��a�Ɨ5.��\�u�-�^�n�LVSE�_[0�Tƶ=�g��
�����hd�Җf�l^M��(�RV�j����R��¨�U�u>��4��<�,�K!pb25��	E @�(�D�'��X=��z�{5�����_������ci����)�X��h���Ͻj�ˢ�;�Y�ly�V�N�1u0vl2�v�^��\�;e���;�4�{
ULz=��$��{Y�T~%�,��l���·�s��Q�ď��=�-�N/垫K�&��N��F���W��g��e�����y���G��h�W߾��g��:d�y��yGN�g�m	�)���7�K����<سG�ݳ�����>��58t�yIx��p��紥<���0���ֲ����)#���&�KLf�Щb�]���3)��-�Lti��ո���׻iY���Y�r9)&"��>M&�V�ے�)�&�>��(��d0�<`�vG�2[��)-;�Q�����JT����;ݔ�G���~��T�B_	&�8G�@��Y߬d�w��:ҝ�_[8r�e�n��'��ő����QP��+�s>����h�[�'����G5
��xЖS잏N��S,=V��U�#���M���������#H<O���Y�ө��,���̥J(���R<�ĩ�w)��$�)�����N�P�3?
���StZ��yV,Y<��݌�7��4V�5����"�k0sz��f����v��d������!^W�+i��/�����*��J��dû�|��˥���M��Rt9NE�����h����^����:��a�>�L\�uV���������w��t�ʤ�b���J��M��QH��C�?�xy�h�=L%�M�jy�Ca�4g(�
���k�3�j���/\�n4z ��ߋ�ɰU�k'���a1��UW�Z����uN�ES��g��bwbt��7L�V�96I�QŷK8X��ɱ��h��90�#76č�0��eGG���t�;Uj��n��V���.N���k����kz�a���?ꟷW�Ú�ƩU���!�8r�����)���~�