BZh91AY&SYq�u� �߀Py���g߰����P (  �RO�4�CF ��4��b��A�ɓ&F�L�L0&&�	�&L�&	���`LM&L�LM2100I !0&��� Q�m@0�6)䟩5_%rDa	�>�U,��Gң�*.�T�)B���ZC
H����T��w�'�N�cs���~��mtJ�_�Ĺ�e��ӻ�J�eYM�/���>Y�Rnmn�5�jX�#+	cbI�6�+�.g��_�^���)^��a�g����\�Z.����tO��Y¡����𞾲�K�C:e_LY��s/\�*Uj�x���'��J*VUUUJ�YQ�;���l�._E�]��MEc���ϥgL%�T/��E�Ti���cQ�k+�Th�t����|:ɹSA�a�������bM!h#X�c���c�N_s��uݔQ�������~Q��;���v��d|��K7i�(�F���O��}F�/�}���^���I6����l�KF�</z�.���a�.9i�ˇ��͏9�WM�oDJ���Գ�]�كL>�cV�}��l_�l�|4�{bR3��t��}����˚+lQؘ���/|c�8G���~RX��I���6��h�q畲�S�y���/�k����b�yS�늇S�����%0��Z�k��5d��k��{���UR���+��a!�J]?�����-�i�:*YS�	4ƈ�bcd]�]s;gokɄ��7�<~�zO��m�7��=�G��3�����Q�^ޣ���=Nx��:9$��T7��a��z8�c�dx��+���uT��<���ÇNx�L���_0]lrؚF�65m�gV��`�b߁B�r9���9Ii.kC����hm׫��ZO遦�&ؿg��R�&�:��֙��"�(H8Һ׀