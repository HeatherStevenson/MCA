BZh91AY&SY���� �߀Ryg���o������`  �     !)�g�h�CC@h �&M4� � dɣ��i�0LM4��8ɓF!���`��i�5S�U)�         2dшbi���4�&&�h �IMd4h1I�
yM`:2AQB�8l?��d���M�& �3����	Ͱ���u��������L������{NX^M_�Z�ED6�YP���C*�.)5]d�ER����Q�]#(�j��--��o�|}�7��n0�-�������<�z�v0ٝ���K�1W>��U�YϞL6i����q���֎�*�j��ȵ�+�ޓ��4a8�V8�5�S5Xsf�u�0�fѷc�������Y��պ�ָZ>ȕ�Tq����H#�~Ll�N�:�wo���z�����m���\���U��:[bnTT)]W�~�ZM�;?��m'V�L��tʲ��2�}i����͔٤���U#5I�BwӾ�J���ch��7}��]O�9թQ��}&&��K�U�4��S���-moW͌M����ՆMk����)�R��%uD@'i�I� `    
h�.��c���=�U�����*�v~�Z�T:������j좬��j{�,��m�ہ�k���9qe�
iFx�:���剥#㢩U,Ѭ�y5��TlP��7UY>�%R�U�ŅTk��Z����P�@D��<�؊ 9�r0�����="c�mv�v��KO�m�v��ɝ���?���Ś)�X������o����c�����e��m�#��f�����5u����:cF������t�?|�|H��B����U	d\{����_���k��D|$�gu���OឫK��g�Q��bt��W����gŞw���y�6��jZL�]�Mc�YD�fl�c{O(�j]��FTb��)��_�v��]�=�c�ɢ?�����{��4���%&$���\Zz{JS(ٽ��J�QoZ��g$�d]�����,�Zg6��7�11=l����C�sN����*��{�9�~�����Gluu�{�α����=�����gj�z�QN�6�B�$u{�FC�������h�l�
KO*)=�iL�y�r�J��f��G����9,�/<8LZ]R��/�8Y��#��Y�3v<���O#'ɒ:���]�O,��7td���l�qP��W�u"�ۣ,{M����'��є�u(�uwr��ʟ\x�7ω��C�kD��j�F�~�Q��|�1$t#ka�tX}���bʋUT���)R�).��#�Z%M��N��vE���go�4��H�i"իStZ��yV�E�S�R[���o߲6+t�/�J��d���1�O���Mv���d�/dnC7��;�?�m�D�n���E�3�rEC�蔠��wLy2�o�7�7:Ⓥ����d����ԼZ*;\�V���5Xx�����ꪴ���:����ܧ7#�ڪOc(��ID�ɪ0(�K�,����cͩ��=,K���$�y����d�J4�D�<�ֻ�d���X�4L�b��=*�l#��Æo�F�Wa�y׏#%�J��ۻ���u��8�:�>M���H�h�1�WJ5������ʏy�0�mF�$q��_�Ͱ�oO)=�����FH�ӮO*���=�����r9%�ê��dvF�q¢���h�-(�n��O׳��إ�U$}��<NN������H�
�]X�