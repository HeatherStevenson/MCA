BZh91AY&SY"M�� ��߀Ryg���o������`1��@ DU�E
(N�@ ���.�*8 `i �w=ފ).-B���7TPIXФ�pYB���ŀ*����j�R`�A$@�&&�M5Q�i��Pz������dh5< R��L�� F� M2` i�I�Ѧ!�A�d�4 ��) �� hh 1 �4  h
R��di�zS�)�4�=OS�P�������Dʥ#I���0!�A�L��4&���*�'�*.�I[U)G�-�G^����M�(��ɥ>}�?��������>���s�c��ҝ
���ܒ��Z6�˷<����EE��|s�}��m/� 2*���HH"�.�/e���C�}�t�! N��'9��y]���>�����]��%�_�|s9���z��w���DI#x�-:�Ch��ɖ�k�a2�ݨw�(��m��5�\��IZ|�st�p�C��F�ȫa��m�ղ>�7Ŷ͘a���_v<�ڡ�Kur�#�Or���C-�nk�r^��gX��ө+��GAg�Iø5ʨi2���j�#�Je����U�v��.�ۛ�n��ڔU�qٗoyh�i���.�'HΫv3kz�E:���7���U\��̬�QV<����m�4���m�7uJ��u}4]F�wb{#���&��.�r�v�kZ��(�b�6�hG��h;�54�iC�E4!�t���G^������]��HSU���ɁS%Ŕ�-��9������أM���F�<}�xI!Y��;�M2���6���5�%��nNA��ڗ���4����q���
U[!Z�������-�:��Db��q�d{4�Y	���2��c��� �����|Kټ�L�h��"Erw||�,7hiV!�M�64�B��P�kz�8t@�M,�rX��t�6��H5��(���x�Ki�$-�2A�z�����x7[牥�l�u#�*䀋#2�9��I=P{w.�H�h�Qvv[�A.w�hդ#��[,|�ۈ���"�$�,�|�ŧ"�
Kvd����D@˸b����j�UJ�ڕz�'w�Cf�<�#[�D�P�pZuR���v�!�X+����ov�\��$k0B:��\J��Ir��1�ݫun��	�Q�H[#54�Xn�UUja�i(H>A(���S�ݏ�r��Ujfٓ �KP�Q
SUvD���$$`�{�&�@��I3X+Sʌ$b�5Zj��U�<�Y��^~ĉ}��c�"s�H5f��HR��AQ�n x�ݹc�S說U�4"hKZf�#��;,���@���Ue7``v-��R�D�N'�Շ�V¤����m �P-j@�qD!V��*�XZ��� I�x B�bz<�Q�d�+E�X��7�*Ʃ+]�y����]ǅ�z�����4���F��+S54�-B��0�@��M
6��
��Q�x�bK\�F!=E.M��&��BmH�Ee��m&�-5kU �Hc�(-���6x��w�.��v���V&�Ey���H�ۛq��ʴ��n�blJJ<i(�L�J�tP�f��,M1 K@�����u=*&[�\��DX���DO ,*�%�+u^ ��`��P�
���7����T*/�TA��d�"���V�U��65��i�B�bm�;��S�Q5���>g��y;��I��_@��d3���j:rJ�M�yJ��{6�U��Ioy���o"	k�1<Oq�ЛǨO\M�	4]�r^�n��F͛k��2T��+�lJͣn=^5ד\��{^ݷ�W�4��"H[��;.I�I��f��^,Wm�x7[�o"^y�yL��jLH$�(��F�ȱ����ZT�W�B a0`o*�H͑����i7:H�u���O/)�J0�o7���m���<q5y��v�����u��]]y�w��)v�h���	o�tȞu�b�z�sH���_V�Y�6!��H�DCW�]����/&���wIn�o�漯b�_7Ƿ����$�"{�yu]��y�Қ��n󉱱����%��3B �ğ�`�.*�eMqn[d2�0n6�7K��ت��H�����!	$�S�t�K@��v��I��������yJ/E�夢�,gOe���Z���_���_��� fa!�
���1P���?w��|�JH�X�Ȕ&�K(��c"�&��c%��E`�X�5%	4��D���
-Ԙ��5)�&���h3̴�Yᖬ�Ql]_����8��?�AV&i��XA^m�^_'ͳ�������٤vy�éؙ�d�B����FQ⎌B���ɓP���^���)W5�Ǉ��Us2���4�Y'0��̷T�	�B��;5ج�=��*���V_<�	[7�z�X����Z�b��J�*lx۵g+3�֤��/`�]x�1w��8X����W:�#���bo�e�]�ٕ����J*�\��s^�S��⼓(�<�R2��eK�R���!u��9ޙ�:ޗ\���nt���������eB�	���,f
���ka����v|7e�ck�}��sk�!�_��80��{ލ}��1e��e�S*�u�!]B��+�{�ہz�2�]������6�l��j�Ab(�ɱ��|u��Z�W�J"�W6LF�I�&��|7������lf�mS%*#jZ�	a���+JH�QH��4�	���J�i�T3b"��
F �1clI d�#J�l�32����R61# ܛ���w���u3э�U��4������L�kѤ�IX�LB��peToN��*T��gbI\�/6��+�Z���c�t;x����i�H����!���G���uiػ&2N�X<i��s�/,2��b_�]W���F�j�)8<tz8�����eaUU�p�e�9k��X&��3�
$ ��_�]��Q$�SY�|����_us��E��{<�����&?��*����e�U%��k���U���{U�=�^Ɣ�����\gl��!o�et��hm�f]��|�c�B�4�����z����ͩ�.���
���ݑ��N��s�HL�e�t�ܬ�����z�0�Ia{��C�o﨩�*��P���}�;��> y�y$T�0�ۋ�b��ѡ�x�B�h�ZJإ!�]�Y�D!B�2�2O��$�S$�.�T�db���bL��[uj�]+s��zm��Ϙ�|k0�HF녫��r����Khn��x� P0M��Lh l4BQoV�5Vb�F#1��&,����k��mk٣Q�I��U�UF��[l&fQ[���aU2ђ���D0�H|��6�.���חh)=:x�D�Ƅ߷��ھ��k%WT�ޱﭯ���n�q�]%���K):�I��@x�Q2��F@�Nqˈ�;*�Rf�(��
�w��a�.��ZY���ý�r��>��1�����Q�*�x��	zZkh���I�)fr!�5'vn���3~T��uB=i��+�P�"	0�@0�
����c�� ޼,�p��P�h�?I��f�OL�vuI�%���;9>|]�Z*]ܗ���z���:98 ��Qx} a�'�"5	�*���o"uX6f�9��V��9{�W�3����QrN�J�^�r�h�����e{��I�9�׈��wq�u��
N뭸���2�Is���6�@�lV�a��k�/�T��#^�����9W �Z��~a� "[��8ix Ðg�������;Ղ���e�y���"YxW{G��h���Cws[�mO�n<�>-��ݿ����d��Į�r�!�·t����ӛ�~�x���/���$�C:d��'�J�֩W�&{�xr �ۇ}����jJN��e]ɽN6��V����~�����Y��V��87��x��7��KЦN/wtpY��� ����W�%�~�B��^�FL�t��MGL�m��4� �K��T�̙-�/��"����"Ԝ⣤qJ �eg����L�!�Җ�i���$4�O  ˾./�ze�2N��X�p��d\/�/������Z*�^�=�.S�V���^j���c$�=�a��p�����������lh�D��\ڄ��%ss�M$�Âg7�t�-Y"�.+<p��E��+4�us�]�u�D]�y�3!s��fq�
���W F�	d$��K
@֖Ф�D�)*_�������d��v�U��RK[�����7!����c{��W}v�n]��͝���EUI8�&&�W��}������z��@��=�mp�[,5n#5��Gn�u�ޫ�eu��8�n�~�H8x��'�R� m�P�N�]w�w*��.�9����,c��-i&*P�Q��������#WU,(�S��v���2
��7���K7ʏtVo�BH�G,��y��w=�m��Ϣ��}����//f�c��՞#�ĝ�����y @؄!���IiD*��I4��3�8���t�x�Z��f,2�8��
�Յ "VA9D�M׈'=�^���d��1����Ղ4aw��`w�{���.�����؈��f& V�\6��g���>�c#�M$���m�ң(1}�����������#��Sd��L ӫ�x�N�VPRk���0ŗ�p�wSm������L�������co���m��`�wu�p�]�1�ҔE9Ѳ D�ws��w;���Qۻ��Eb�V7˕��5�ZѠ�F���E�,T�EQ���Q�[Ɗ�EE�����ڍLm�o���uA}#O��8��U`�`�}�� ��a�������� Z���2	Rn�x�
�'f˨���]{��Zk�7���	�>^�υ����T�ޱ��� :x�;̕�o�o�,hI4K,=���&�2��}+���uB��3��d���/|%��g�|9$�*�b�|�|�R�*�c��&���:�F6�;i�<�T���dyB���n�M�Q� �pvw��A�4�^NY�!uy�b���߮b��s^���Uy\�r�=�QG�a���"2�����f��m5�ܳCv��vŹ8q9-��ٝG%�C���/�?X���H I����*(���wi4�tN�W{�1��қ53PJ�UJ� �$8p?S��߷�w��t����Og�2��
�Z^�#�'0Z�A6��M���)���-�ם]F���|���D��Ѩ�A������04�a�`�E
I��X�f(�b�T ldѢ"iR�`��
�	i���" ��Ld�-���B�ƚm�H��iJBK�+YF{G���Vw�bA�ϫ�b)�����K2�qqM��,,����{}d��uYc�VJ	)vF�yW:��W)L�g��3τ�i>0�y��E�$�5�1��,�5qt�B�qO&�����+BߨUZ��r0PnK*��̩���m�o7���i��6�őkN,X����w-�'�TL����1Q�=�ݤVb��FkP�A�����ϵ})K�s���j�ٸ��ғ�M�gA)I��Kjn�*��7%g���y�:\�#��p ��%T[��rI�n����*��3����QHC��sg;�9���JY�I��ܜ�#e�r"�f�����HF�L��|<\��٪0,�[�I^͒�3��5��L������}�{A
��þ��|��F�QV,Wü}���!IC�6)rV-����b��BM(��\����.�n򾲬�m�(�`�i��*%fɡ4i
��R4�A�I5mz�}T[cl ��k��V�yK9��������Ҳ��bH�6	�E �P�in�W�s���Y�����8�7��`��ꔵ��X���$��&c8z�Z=��`y���ׇ�N�=��� Ik4�߰Ȋ�ˊi{n
\<E�I�eb�0���{;B@�ȿ;�绲;��f�~骏(<�����uTpkT¢�!a>�����w�kk8t��C��"&;�*
���OX�s�y_��b����%!�8�6��9���R�1B]\�O��a2Q#1DɄ�=�/���PA��_���@�x���<B���!	���;���@kHm	��@������%�Z�4f���-���w���>"�/<��z�m�bR��$�Q��j6��hDh�˛�b�.s��F4�D&�}�6D�bw|�6��O��E�'V+�����#Nњ�)^���4a	X�5w�Vx�[E�ʾ���ˇ �j���uV;��3�B���˕x�}A��8�!�B@�;�&ġh������y�cΗ�Wi A�\�)b���9��Ҏ+]'����&����T{��l�%F��vA�K���  ��	�F��,��4�+6'�ɺ�p画�V�<�sOZ��$��6c��1b�H8iA�wѾ�ja����r9$����y'��*���m������KOI����ⱍ��5}�h�UuWu�4�}��BKl<�z�3Q��O�H��������F���#1qt�T�=�S'b:���X�FSF�ҩp�ӥ�`���GoA�S�g�$�%��;����� �8[)C��]�*O'z����"�2X1E�i�|����F,d��l����������qG���l���*�N��(�#Af��W��f<���w��"�#o�pۛ۷|r����v��'3�����T�BIBHq��SzѦZ+�m6�R���[ڸgW9�{�j�kO��Η}���a����WL��3"]U�'n�}v��O7����_]��=�q+[��u<Z���W���7���1���ܢ�"��4�Z���`���^��}��O��eE-��\+���>�_��:��L��/HHXcӊW�L!��͊/8nhP$��H��d��%xtC�R��7ڨq^Z���W�co.���s�Y9S�/���?t��r����Ɍ�[m��6�]Q��ݜz�5��
�2�:O."<��m�\��BTJ��ۼ[>��>߷h���6U��!0+��!9���G�25Ư��!�,rsV���k�٘�h��l�{�-]@�I����5b�x1���u2ڢNzN^x�gzfaw���7����P���%�=�נT�'���q߫�1��w�j30��336a�(�f��ڒ���4l��rpm٣��چ��Bճ��88%omr��=v�6����[3jX�+LL��&��i6e3mh����սƶ��{4�l&FUVF#%��c�,���a!�"��i2�L�aMD42bə*� hda�,Ča@a�$ʈ`�@	"Zl*�af1�
FX�,=+����� m	��߈]�������,�7|�Y�"�;��C�����x�RV_��9��+4���^X���pk�5f��ƵL�
�qIP��L��/Xn6�y:������I(�
Q}�]46�����?�ɾ\ۏa��і�����Zy^c����WO�%/w'Vl>�����:��ţ�#W9D�&�uR(;4,]���RLJ2Q��V2��$���b.V<PF�ݍN2J��$ �L��aX�0����I��6��b2K)1UeFJ�Q�dF(�ʦ)d,I2)eLQ��K$`�	�#�X���L*ɒc	�*��U�֥��.���\�Zxa��\�>����IEťj��#�/8��E�6��a7�yu��c߈T#ݯӣ�u�̒���ǭlu�NMi)@��N���+�f�-Vǒ�*���d,QZ�x�s���U��Ԉ��>;�t!�_v��W���ܒ�^b�2R���L�v����Vi���1�ŷ��V�*-�)(�-�~!��u�aױ��=C�J.f�m�p`�7/[�JJ/4�u��Z�����EIbL<y��!���O��H!�9c�0ZE�����NSM�?��y��eBh�QcL��84�~�O�Y���t�RQ}&���:�.��$��{�q�k��q�k��8u���nƌyNw���c�p��á��z������(��̝}���G�����w����nY���㡜�5�E�B`u��,��2t�N��C�|�2��DS�(����)���B�@n�6L�x=�q�p�$
��'pw��2ѕF� �㲗�гr-aH��+&:83V3:A��!a,=��	��(�����z�'+]m%{;�����-Ɔk��B2-��8Y#/b�J��i�o�a�����f�s��.�p� D�/h