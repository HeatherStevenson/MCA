BZh91AY&SY�Ny� �߀Py���g߰?���P��*�@�IB�bDcA0����#Mc�2b`b0#L1&L0H�2�M54�6��   H= 挘� ���F	� �D&�i�bS��jbzi22 d�d� �k  �H��Ͳ Y2�.P��!�H!}�"B'|%�F�8Bxv�T��&��O�(�xCXl��Hj�U����pa�A^�4��� �fL%d`;�%��SITv�Z� �4���m�{L�s�Ʈ@]0)i�;�/�B��e)	ܒ[)�q���~-a�2��!z��ԩ,�����[ʦ4ә��m�@��X� �1�0��I*���N�l�0U�!�d��a�Qx�U	�)9�*jf�b)es���y�pxO�G��ӡ�wI�H�F��q3��'�~��n��R����M�K4�6��5;�F�c�XE�L��(6��MX���̑��8?����_�E�(3���|u}ع@R����\B��0m��4y�_O_�ȿ|�a)U��$WY&k�Z��=�`Pٔ@�Z$�[��xGL݁���f�A��4<�sذh�y�"��=�ޔ�F��	�t<=�CP��������8x��Ǣ�0,�A�9$Ѥy����\�+�lN�u�qP�d 쩴��H��FU�1�����G�3�0�꣊]*��)ؐD�J���+�;�R�pN�p�!QZi�`X '*|��-�\"��B�lXDʅa�܎���R ��΃������t�7
&Mh�?GU)F����ގ�9\�2�S�V�'�C���׺s�ug�lu�z�e� e�b�ޱ�Ʀb.��#�(nٽ�������)k��힔�"� �f7�w$S�	�p