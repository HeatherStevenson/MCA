BZh91AY&SYq��� �_�Py���g߰����P��j
�$�?U�MM<�4�A�d� 4� ڃ�A�ɓ&F�L�L4�����4�� Cё�h ���a2dɑ��4�# C �!MM�jyM�@��S� M4fI��8"���A#P}�H`)C�B���Z=0�a@�	Ո�t��
���$����6�5��e&��y��3$�j�GƸ1��'�3��k|��iY���Q�1Ĉ��?s��]� ���Y.	��u0k��H�Y��0����T���2|!���I��Mk���ZS��pȪ��=Q�طd�jAU	ADD@{z�q�h�+(Ĳ�Sb_L�3D���A�:P�"�
\��r�6C"F�f���,�")���*O���륎�^�&��$|O_��=8h�쓚������½�҇*��\S���n��-�7ɳ���$�M�e?>So�@k܁_����򈪑�m�1������R��quf���4m6I���y�!�HH�$�1-)�T�P��c��$Ȯ���^�a�1ַ;�<�N�-Ȱf	p��O�<S-�P�m.M���S	 �
�R6hQ++��(�$d�\,T� ��<����������[A�7��MC qNJ��� :(<(���U��tG�i�:!�HvU4�����N���&��P�:��*,l����n��ό��JԀcPsە���(Xd��Qu]e� �5���Â�BD���G����9Q�(��0%����Mcih^�R�`D�T"\A�DMI�a�����|��f67�v1P�p���_��dh\!Ϩ��J��w2?�bS$��_��1@��4���.�p� ����