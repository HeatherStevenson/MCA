BZh91AY&SY���� �_�Py���g߰����P��T(�$ښG�2&OP�i��� � 挘� ���F	� �j����h4�  @ 9�&& &#4���d�#Q@ji�d�i5=�bh�'���EF� �
`��� ��=��)�`+C�B�.�^<Жa@����CW�8Md��P8F؆
�n��$�yz��7D��I9Pu�t:���c<�u�3���:�@0�GRg�DnJw�N�,�<� ,�	�l���z����IMQ�����7BZ� ���@*d;��Pm3BO01!�<��
�I12@{�'a��B�Ђ��%�C���,|Lf���z�����������W��!
&ɱgH��)��w?���(�r#䳡�O�T��-�>�ݹdAb��ENp��J�w@��������%�I�h�qZ'������zA��	5�\ZY�*�ȳ��~Q�c JY=�;�)Nr�=\���-3B����_y�N���Q�
@�Et]�i��}�����Nv�I�]��i.���#G0݃�h}�pҰdR��:J�����t�G3K�����y(�TL+�����gP�+�7T�XY�=) l�<���A���rober-��*�@⟎��� 9Px�#E�2(�z��G�i�8C��9��v�i4M8���<)QcnA��4јu:����5�e,Q�
���zs+����R˔@��0���ԑ q8r$|>g�u�����G�����F�6lߍ��7�lRo��̙�n�NTۨ�k�lu�4����yPֿ��dhk��`SyC�>�{#�x`L���fɈ"���n���H�
���